module blinky #(parameter clk_freq_hz = 0)
