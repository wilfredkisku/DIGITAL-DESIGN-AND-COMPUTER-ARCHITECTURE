module encoder32_5(en, A, Y);
        input en;
        input [31:0] A;
        output reg [4:0] Y;

endmodule

